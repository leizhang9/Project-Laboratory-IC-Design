----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 23.06.2022 11:04:11
-- Design Name: 
-- Module Name: tb_modify - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity tb_modify is
--  Port ( );
end tb_modify;

architecture Behavioral of tb_modify is
    component modify
        Port ( clk : in std_logic;
           fsm_alarm : in STD_LOGIC;
           key_enable : in STD_LOGIC;
           key_p_m : in STD_LOGIC;
           rst : in STD_LOGIC;
           ss : out STD_LOGIC_VECTOR (5 downto 0);
           mm : out STD_LOGIC_VECTOR (5 downto 0);
           hh : out STD_LOGIC_VECTOR (4 downto 0));
    end component;
    
    signal key_enable, key_p_m, rst, clk, fsm_alarm: std_logic := '0';
    signal ss : STD_LOGIC_VECTOR (5 downto 0);
    signal mm : STD_LOGIC_VECTOR (5 downto 0);
    signal hh : STD_LOGIC_VECTOR (4 downto 0);
    constant clk_period: time := 10 ns;
begin
    uut: modify port map (clk => clk, fsm_alarm => fsm_alarm, key_enable => key_enable, key_p_m => key_p_m, rst => rst, ss => ss, mm => mm, hh => hh);
    clock: process
    begin
        clk <= '0';
        wait for clk_period/2;
        clk <= '1';
        wait for clk_period/2;
    end process clock;
    process
    begin 
    wait for 100ns;
    key_enable <= '1';
    key_p_m <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    fsm_alarm <= '1';
    wait for 10 ns;
    key_enable <= '0';
    rst <= '1';
    wait for 10 ns;
    rst <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
        wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
        wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
        wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
        wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait for 100ns;
    key_enable <= '1';
    wait for 10 ns;
    key_enable <= '0';
    wait;
    end process;

end Behavioral;
